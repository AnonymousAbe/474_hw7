module clock(
	input			reset_n,		//reset pin
	input			clk_1sec,		//1 sec clock
	input			clk_1ms,		//1 mili sec clock
	input			mil_time,		//mil time pin
	output reg [6:0]	segment_data,		//output 7 seg data
	output reg [2:0]	digit_select		//digit select
);








endmodule
